-------------------------------------------------------------------------
-- Colton Hazlett
-- Department of Electrical and Computer Engineering
-- Iowa State University
-------------------------------------------------------------------------
-- tb_dmem.vhd
-------------------------------------------------------------------------
-- DESCRIPTION: This file contains a testbench for the ram
--              
-- 01/03/2020 by H3::Design created.
-------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_textio.all;  -- For logic types I/O
library std;
use std.env.all;                -- For hierarchical/external signals
use std.textio.all;             -- For basic I/O

-- Usually name your testbench similar to below for clarity tb_<name>
-- TODO: change all instances of tb_TPU_MV_Element to reflect the new testbench.
entity tb_dmem is
  generic(gCLK_HPER   : time := 10 ns);   -- Generic for half of the clock cycle period
end tb_dmem;

architecture mixed of tb_dmem is

-- Define the total clock period time
constant cCLK_PER  : time := gCLK_HPER * 2;

-- We will be instantiating our design under test (DUT), so we need to specify its
-- component interface.
-- TODO: change component declaration as needed.
component mem is
  port( clk		: in std_logic;
	addr	        : in std_logic_vector(9 downto 0);
	data	        : in std_logic_vector(31 downto 0);
	we		: in std_logic := '1';
	q		: out std_logic_vector(31 downto 0));
end component;

-- Create signals for all of the inputs and outputs of the file that you are testing
-- := '0' or := (others => '0') just make all the signals start at an initial value of zero
signal CLK, reset : std_logic := '0';

-- TODO: change input and output signals as needed.
signal s_addr      : std_logic_vector(9 downto 0);
signal s_we        : std_logic;
signal s_data      : std_logic_vector(31 downto 0);
signal s_Q         : std_logic_vector(31 downto 0);

begin

  -- TODO: Actually instantiate the component to test and wire all signals to the corresponding
  -- input or output. Note that DUT0 is just the name of the instance that can be seen 
  -- during simulation. What follows DUT0 is the entity name that will be used to find
  -- the appropriate library component during simulation loading.
  dmem: mem
  port map( clk  => CLK,
            addr => s_addr, 
            data => s_data,
            we   => s_we,
            q    => s_Q);

  --You can also do the above port map in one line using the below format: http://www.ics.uci.edu/~jmoorkan/vhdlref/compinst.html

  
  --This first process is to setup the clock for the test bench
  P_CLK: process
  begin
    CLK <= '1';         -- clock starts at 1
    wait for gCLK_HPER; -- after half a cycle
    CLK <= '0';         -- clock becomes a 0 (negative edge)
    wait for gCLK_HPER; -- after half a cycle, process begins evaluation again
  end process;

  -- This process resets the sequential components of the design.
  -- It is held to be 1 across both the negative and positive edges of the clock
  -- so it works regardless of whether the design uses synchronous (pos or neg edge)
  -- or asynchronous resets.
  P_RST: process
  begin
  	reset <= '0';   
    wait for gCLK_HPER/2;
	reset <= '1';
    wait for gCLK_HPER*2;
	reset <= '0';
	wait;
  end process;  
  
  -- Assign inputs for each test case.
  -- TODO: add test cases as needed.
  P_TEST_CASES: process
  begin
    wait for gCLK_HPER/2; -- for waveform clarity, I prefer not to change inputs on clk edges

    --------------------------------------------------------
    -- Step 1 is transfer the data from memory 0x0 to 0x100
    --------------------------------------------------------

    --Transfer 1:
    -- Read the data value at index 0 and store at index 0x100
    s_we <= '0';
    s_addr <= "0000000000"; --Reads value 0
    wait for gCLK_HPER*2;
    s_data <= s_Q;          --Set data to the value that was read
    s_addr <= "0100000000"; --Write value at index 0x100
    s_we   <= '1';          --Write enable 1 tpo activate the write
    wait for gCLK_HPER*2;
    wait for gCLK_HPER*2;

    --Transfer 2:
    -- Read the data value at index 1 and store at index 0x101
    s_we <= '0';
    s_addr <= "0000000001"; --Reads value 1
    wait for gCLK_HPER*2;
    s_data <= s_Q;          --Set data to the value that was read
    s_addr <= "0100000001"; --Write value at index 0x101
    s_we   <= '1';          --Write enable 1 tpo activate the write
    wait for gCLK_HPER*2;
    wait for gCLK_HPER*2;

    --Transfer 3:
    -- Read the data value at index 2 and store at index 0x102
    s_we <= '0';
    s_addr <= "0000000010"; --Reads value 2
    wait for gCLK_HPER*2;
    s_data <= s_Q;          --Set data to the value that was read
    s_addr <= "0100000010"; --Write value at index 0x102
    s_we   <= '1';          --Write enable 1 tpo activate the write
    wait for gCLK_HPER*2;
    wait for gCLK_HPER*2;

    --Transfer 4:
    -- Read the data value at index 3 and store at index 0x103
    s_we <= '0';
    s_addr <= "0000000011"; --Reads value 3
    wait for gCLK_HPER*2;
    s_data <= s_Q;          --Set data to the value that was read
    s_addr <= "0100000011"; --Write value at index 0x103
    s_we   <= '1';          --Write enable 1 tpo activate the write
    wait for gCLK_HPER*2;
    wait for gCLK_HPER*2;

    --Transfer 5:
    -- Read the data value at index 4 and store at index 0x104
    s_we <= '0';
    s_addr <= "0000000100"; --Reads value 4
    wait for gCLK_HPER*2;
    s_data <= s_Q;          --Set data to the value that was read
    s_addr <= "0100000100"; --Write value at index 0x104
    s_we   <= '1';          --Write enable 1 tpo activate the write
    wait for gCLK_HPER*2;
    wait for gCLK_HPER*2;

    --Transfer 6:
    -- Read the data value at index 5 and store at index 0x105
    s_we <= '0';
    s_addr <= "0000000101"; --Reads value 5
    wait for gCLK_HPER*2;
    s_data <= s_Q;          --Set data to the value that was read
    s_addr <= "0100000101"; --Write value at index 0x105
    s_we   <= '1';          --Write enable 1 tpo activate the write
    wait for gCLK_HPER*2;
    wait for gCLK_HPER*2;

    --Transfer 7:
    -- Read the data value at index 6 and store at index 0x106
    s_we <= '0';
    s_addr <= "0000000110"; --Reads value 6
    wait for gCLK_HPER*2;
    s_data <= s_Q;          --Set data to the value that was read
    s_addr <= "0100000110"; --Write value at index 0x106
    s_we   <= '1';          --Write enable 1 tpo activate the write
    wait for gCLK_HPER*2;
    wait for gCLK_HPER*2;

    --Transfer 8:
    -- Read the data value at index 7 and store at index 0x107
    s_we <= '0';
    s_addr <= "0000000111"; --Reads value 7
    wait for gCLK_HPER*2;
    s_data <= s_Q;          --Set data to the value that was read
    s_addr <= "0100000111"; --Write value at index 0x107
    s_we   <= '1';          --Write enable 1 tpo activate the write
    wait for gCLK_HPER*2;
    wait for gCLK_HPER*2;

    --Transfer 9:
    -- Read the data value at index 8 and store at index 0x108
    s_we <= '0';
    s_addr <= "0000001000"; --Reads value 8
    wait for gCLK_HPER*2;
    s_data <= s_Q;          --Set data to the value that was read
    s_addr <= "0100001000"; --Write value at index 0x108
    s_we   <= '1';          --Write enable 1 tpo activate the write
    wait for gCLK_HPER*2;
    wait for gCLK_HPER*2;

    ----------------------------------------------------------------------------
    -- Step 2 is to Re-read all the data to make sure it transferred correctly
    ----------------------------------------------------------------------------
    
    --Read 1:
    s_we   <= '0';
    s_addr <= "0100000000";
    wait for gCLK_HPER*2;
    -- Expect: s_Q = 0xFFFFFFFF (-1)

    --Read 2:
    s_addr <= "0100000001";
    wait for gCLK_HPER*2;
    -- Expect: s_Q = 0xFFFFFFFE (-2)

    --Read 3:
    s_addr <= "0100000010";
    wait for gCLK_HPER*2;
    -- Expect: s_Q = 0xFFFFFFFD (-3)

    --Read 4:
    s_addr <= "0100000011";
    wait for gCLK_HPER*2;
    -- Expect: s_Q = 0xFFFFFFFC (-4)

    --Read 5:
    s_addr <= "0100000100";
    wait for gCLK_HPER*2;
    -- Expect: s_Q = 0xFFFFFFFB (-5)

    --Read 6:
    s_addr <= "0100000101";
    wait for gCLK_HPER*2;
    -- Expect: s_Q = 0xFFFFFFFA (-6)

    --Read 7:
    s_addr <= "0100000110";
    wait for gCLK_HPER*2;
    -- Expect: s_Q = 0xFFFFFFF9 (-7)

    --Read 8:
    s_addr <= "0100000111";
    wait for gCLK_HPER*2;
    -- Expect: s_Q = 0xFFFFFFF8 (-8)

    --Read 9:
    s_addr <= "0100001000";
    wait for gCLK_HPER*2;
    -- Expect: s_Q = 0xFFFFFFF7 (-9)

    -- TODO: add test cases as needed (at least 3 more for this lab)
  end process;

end mixed;