-------------------------------------------------------------------------
-- Colton Hazlett
-- Department of Electrical and Computer Engineering
-- Iowa State University
-------------------------------------------------------------------------
-- tb_control.vhd
-------------------------------------------------------------------------
-- DESCRIPTION: This file contains a testbench for the register N-Bits wide
--              
-- 01/03/2020 by H3::Design created.
-------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_textio.all;  -- For logic types I/O
library std;
use std.env.all;                -- For hierarchical/external signals
use std.textio.all;             -- For basic I/O

-- Usually name your testbench similar to below for clarity tb_<name>
-- TODO: change all instances of tb_TPU_MV_Element to reflect the new testbench.
entity tb_control is
  generic(gCLK_HPER   : time := 10 ns);   -- Generic for half of the clock cycle period
end tb_control;

architecture mixed of tb_control is

-- Define the total clock period time
constant cCLK_PER  : time := gCLK_HPER * 2;

-- We will be instantiating our design under test (DUT), so we need to specify its
-- component interface.
-- TODO: change component declaration as needed.
component control is
  port(instruction  : in  std_logic_vector(5 downto 0);
       RegDst       : out std_logic;
       jump         : out std_logic;
       branch       : out std_logic;
       MemWR        : out std_logic;
       MemtoReg     : out std_logic;
       ALUSrc       : out std_logic;
       RegWE        : out std_logic;
       immSigned    : out std_logic;
       equals       : out std_logic;
       ALUop        : out std_logic_vector(3 downto 0));
end component;

-- Create signals for all of the inputs and outputs of the file that you are testing
-- := '0' or := (others => '0') just make all the signals start at an initial value of zero
signal CLK, reset : std_logic := '0';

-- TODO: change input and output signals as needed.
signal s_ins      : std_logic_vector(5 downto 0);
signal s_ALUop    : std_logic_vector(3 downto 0);
signal s_regDst, s_jump, s_branch, s_memWR, s_MemtoReg, s_ALUSrc, s_RegWE, s_immSigned, s_equals : std_logic;

begin

  -- TODO: Actually instantiate the component to test and wire all signals to the corresponding
  -- input or output. Note that DUT0 is just the name of the instance that can be seen 
  -- during simulation. What follows DUT0 is the entity name that will be used to find
  -- the appropriate library component during simulation loading.
  DUT0: control
  port map( instruction => s_ins,
            RegDst      => s_regDst,
            jump        => s_jump,
            branch      => s_branch,
            MemWR       => s_memWR,
            MemtoReg    => s_MemtoReg,
            ALUSrc      => s_ALUSrc,
            RegWE       => s_RegWE,
            immSigned   => s_immSigned,
            equals      => s_equals,
            ALUop       => s_ALUop);
  --You can also do the above port map in one line using the below format: http://www.ics.uci.edu/~jmoorkan/vhdlref/compinst.html

  
  --This first process is to setup the clock for the test bench
  P_CLK: process
  begin
    CLK <= '1';         -- clock starts at 1
    wait for gCLK_HPER; -- after half a cycle
    CLK <= '0';         -- clock becomes a 0 (negative edge)
    wait for gCLK_HPER; -- after half a cycle, process begins evaluation again
  end process;

  -- This process resets the sequential components of the design.
  -- It is held to be 1 across both the negative and positive edges of the clock
  -- so it works regardless of whether the design uses synchronous (pos or neg edge)
  -- or asynchronous resets.
  P_RST: process
  begin
  	reset <= '0';   
    wait for gCLK_HPER/2;
	reset <= '1';
    wait for gCLK_HPER*2;
	reset <= '0';
	wait;
  end process;  
  
  -- Assign inputs for each test case.
  -- TODO: add test cases as needed.
  P_TEST_CASES: process
  begin
    wait for gCLK_HPER*2;
    wait for gCLK_HPER/2; -- for waveform clarity, I prefer not to change inputs on clk edges
    
    -- Test Case 1: 
    -- Set to a R-Type instruction
    s_ins <= "000000";
    wait for gCLK_HPER*2;
    -- Expected output 
    --    ALUop     -> 0x0
    --    ALUSrc    -> 0
    --    MemtoReg  -> 0
    --    MemWR     -> 0
    --    RegWE     -> 1
    --    RegDst    -> 1
    --    immSigned -> 0
    --    jump      -> 0
    --    branch    -> 0

    -- Test Case 2: 
    -- Set to addi
    s_ins <= "001000";
    wait for gCLK_HPER*2;
    -- Expected output 
    --    ALUop     -> 0x1
    --    ALUSrc    -> 1
    --    MemtoReg  -> 0
    --    MemWR     -> 0
    --    RegWE     -> 1
    --    RegDst    -> 0
    --    immSigned -> 1
    --    jump      -> 0
    --    branch    -> 0


    -- Test Case 3: 
    -- Set to addiu
    s_ins <= "001001";
    wait for gCLK_HPER*2;
    -- Expected output 
    --    ALUop     -> 0x2
    --    ALUSrc    -> 1
    --    MemtoReg  -> 0
    --    MemWR     -> 0
    --    RegWE     -> 1
    --    RegDst    -> 0
    --    immSigned -> 1
    --    jump      -> 0
    --    branch    -> 0
    

    -- Test Case 4: 
    -- Set to andi
    s_ins <= "001100";
    wait for gCLK_HPER*2;
    -- Expected output 
    --    ALUop     -> 0x6
    --    ALUSrc    -> 1
    --    MemtoReg  -> 0
    --    MemWR     -> 0
    --    RegWE     -> 1
    --    RegDst    -> 0
    --    immSigned -> 1
    --    jump      -> 0
    --    branch    -> 0


    -- Test Case 5: 
    -- Set to lui
    s_ins <= "001111";
    wait for gCLK_HPER*2;
    -- Expected output 
    --    ALUop     -> 0x5
    --    ALUSrc    -> 1
    --    MemtoReg  -> 0
    --    MemWR     -> 0
    --    RegWE     -> 1
    --    RegDst    -> 0
    --    immSigned -> 0
    --    jump      -> 0
    --    branch    -> 0


    -- Test Case 6: 
    -- Set to lw
    s_ins <= "100011";
    wait for gCLK_HPER*2;
    -- Expected output 
    --    ALUop     -> 0xA
    --    ALUSrc    -> 1
    --    MemtoReg  -> 1
    --    MemWR     -> 1
    --    RegWE     -> 1
    --    RegDst    -> 0
    --    immSigned -> 1
    --    jump      -> 0
    --    branch    -> 0


    -- Test Case 7: 
    -- Set to xori
    s_ins <= "001110";
    wait for gCLK_HPER*2;
    -- Expected output 
    --    ALUop     -> 0x8
    --    ALUSrc    -> 1
    --    MemtoReg  -> 0
    --    MemWR     -> 0
    --    RegWE     -> 1
    --    RegDst    -> 0
    --    immSigned -> 0
    --    jump      -> 0
    --    branch    -> 0


    -- Test Case 8: 
    -- Set to ori
    s_ins <= "001101";
    wait for gCLK_HPER*2;
    -- Expected output 
    --    ALUop     -> 0x7
    --    ALUSrc    -> 1
    --    MemtoReg  -> 0
    --    MemWR     -> 0
    --    RegWE     -> 1
    --    RegDst    -> 0
    --    immSigned -> 0
    --    jump      -> 0
    --    branch    -> 0


    -- Test Case 9: 
    -- Set to slti
    s_ins <= "001010";
    wait for gCLK_HPER*2;
    -- Expected output 
    --    ALUop     -> 0x9
    --    ALUSrc    -> 1
    --    MemtoReg  -> 0
    --    MemWR     -> 0
    --    RegWE     -> 1
    --    RegDst    -> 0
    --    immSigned -> 1
    --    jump      -> 0
    --    branch    -> 0


    -- Test Case 10: 
    -- Set to sw
    s_ins <= "101011";
    wait for gCLK_HPER*2;
    -- Expected output 
    --    ALUop     -> 0xB
    --    ALUSrc    -> 1
    --    MemtoReg  -> 1
    --    MemWR     -> 1
    --    RegWE     -> 0
    --    RegDst    -> 0
    --    immSigned -> 1
    --    jump      -> 0
    --    branch    -> 0


    -- Test Case 11: 
    -- Set to beq
    s_ins <= "000100";
    wait for gCLK_HPER*2;
    -- Expected output 
    --    ALUop     -> 0xC
    --    ALUSrc    -> 1
    --    MemtoReg  -> 0
    --    MemWR     -> 0
    --    RegWE     -> 1
    --    RegDst    -> 0
    --    immSigned -> 0
    --    jump      -> 0
    --    branch    -> 0


    -- Test Case 12: 
    -- Set to bne
    s_ins <= "000101";
    wait for gCLK_HPER*2;
    -- Expected output 
    --    ALUop     -> 0xD
    --    ALUSrc    -> 1
    --    MemtoReg  -> 0
    --    MemWR     -> 0
    --    RegWE     -> 1
    --    RegDst    -> 0
    --    immSigned -> 0
    --    jump      -> 0
    --    branch    -> 0


    -- Test Case 13: 
    -- Set to j
    s_ins <= "000010";
    wait for gCLK_HPER*2;
    -- Expected output 
    --    ALUop     -> 0x0
    --    ALUSrc    -> 0
    --    MemtoReg  -> 0
    --    MemWR     -> 0
    --    RegWE     -> 0
    --    RegDst    -> 0
    --    immSigned -> 0
    --    jump      -> 1
    --    branch    -> 0


    -- Test Case 14: 
    -- Set to jal
    s_ins <= "000011";
    wait for gCLK_HPER*2;
    -- Expected output 
    --    ALUop     -> 0x1
    --    ALUSrc    -> 0
    --    MemtoReg  -> 0
    --    MemWR     -> 0
    --    RegWE     -> 0
    --    RegDst    -> 0
    --    immSigned -> 0
    --    jump      -> 1
    --    branch    -> 0

    -- TODO: add test cases as needed (at least 3 more for this lab)
  end process;

end mixed;