-------------------------------------------------------------------------
-- Colton Hazlett
-- Department of Electrical and Computer Engineering
-- Iowa State University
-------------------------------------------------------------------------


-- ALU.vhd
-------------------------------------------------------------------------
-- DESCRIPTION: This file contains an implementation of an Ones complementor 
-- that will negate each bit given in the single input.
--
--
-- NOTES:
-- 2/4/2020 by H3::Created.
-------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

entity ALU is
  port(i_A     : in  std_logic_vector(31 downto 0);
       i_B     : in  std_logic_vector(31 downto 0);
       ALUop   : in  std_logic_vector(3 downto 0);
       o_Carry : out std_logic;
       o_Ovf   : out std_logic;
       o_Zero  : out std_logic;
       o_Q     : out std_logic_vector(31 downto 0));


end ALU;

architecture structural of ALU is

   ------------------------------------------
   -- Step 1: Instantiate all the components
   ------------------------------------------
   component add_sub_N
     port( i_C         :  in std_logic;
           i_nAdd_Sub  :  in std_logic;
           i_A         :  in std_logic_vector(N-1 downto 0);
           i_B         :  in std_logic_vector(N-1 downto 0);
           o_S         : out std_logic_vector(N-1 downto 0);
           o_C         : out std_logic);
   end component;

   component barrel_shift
     port(i_Data 	: in std_logic_vector(31 downto 0);
	  i_left 	: in std_logic;                     --1 for left and 0 for right 
	  i_logic	: in std_logic;                     --1 for logic (unsigned) and 0 for arithmetic (signed)
	  i_shift	: in std_logic_vector(4 downto 0);  --shift amount
	  o_Data	: out std_logic_vector(31 downto 0));
   end component;

   component c_gates_N
     port(i_A   : in  std_logic_vector(N-1 downto 0);
          i_B   : in  std_logic_vector(N-1 downto 0);
          i_Sel : in  std_logic_vector(1 downto 0);         --Chooses between and, or, xor, & nor
          o_Q   : out std_logic_vector(N-1 downto 0));
   end component;

   component mux2t1_N
     port(i_S          : in std_logic;
          i_D0         : in std_logic_vector(N-1 downto 0);
          i_D1         : in std_logic_vector(N-1 downto 0);
          o_OA         : out std_logic_vector(N-1 downto 0));
   end component;

   ---------------------------------------------------
   --Step 2: Create all the signals that we will need
   ---------------------------------------------------


begin

  ---------------------------------------------
  --Step 3: Map all the inner componets to run
  ---------------------------------------------

end structural;